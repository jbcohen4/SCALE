Title: AD590 / OutputCurrent (A)
*************************************

*Voltage Source
VIN 2 0 DC 0V
VOUT 20 0 0

*Circuit Core
R7 20 0 1m

*Input
.dc VIN 0 30 1

*Output
.print dc format=noindex file=tempfiles\xyce_output\xoutput_73.out
+ V(2)
+ I(VOUT)

*Diode: D<name> <anode node (+)> <cathode node (-)> <model name> [area value]
**********************************
*PNP
D1 4 8 DMODPNP 1.6 temp=25
D2 4 8 DMODPNP 1.6 temp=25
D3 4 8 DMODPNP 1.6 temp=25
D4 4 8 DMODPNP 1.6 temp=25
D5 3 8 DMODPNP 1.6 temp=25
D6 2 7 DMODPNP 1.6 temp=25
*NPN
D7 6 11 DMODNPN 4 temp=25
D8 1 11 DMODNPN 4 temp=25
D9 5 15 DMODNPN 32 temp=25
D10 5 12 DMODNPN 4 temp=25
D11 5 12 DMODNPN 4 temp=25

*Capacitance: C<name> <+ node> <- node> [model name] <value> + [IC=<initial value>]
c1 1 8 26p

*Resistance: R<name> <+ node> <- node> [model name] <value>
r1 2 4 260
r2 2 3 1040
r3 5 16 5000
r4 11 5 11000
r5 12 20 146
r6 15 20 820

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q1 6 8 4 QLPMOD 1.6 temp=25
Q2 6 8 4 QLPMOD 1.6 temp=25
Q3 1 8 4 QLPMOD 1.6 temp=25
Q4 1 8 4 QLPMOD 1.6 temp=25
Q5 8 8 3 QLPMOD 1.6 temp=25
Q6 7 7 2 QLPMOD 1.6 temp=25
Q7 7 6 11 QNMOD 4 temp=25
Q8 8 1 11 QNMOD 4 temp=25
Q9 6 5 15 QNMOD 32 temp=25
Q10 5 5 12 QNMOD 4 temp=25
Q11 1 5 12 QNMOD 4 temp=25

*Q9, Q10, and Q11 emitter area still need to be cal

*JFET: J<name> <drain> <gate> <source> <model name> [area value]
J1 8 16 11 NJF_TYP

*Library
* npn prerad off ctp 3b
.model QNMOD NPN (              
+IS=2.354912E-16
+BF=84.058
+NF=0.986787     
+VAF=351.9861415
+IKF=9.86E-3
+NK=0.47574  
+ISE=7.1029E-15
+NE=2.06453  
+BR=0.697       
+NR=2
+VAR=100
+IKR=0.1         
+ISC=1E-17
+NC=2                          
+RB=140.86       
+IRB=1E-3 
+RBM=50                        
+RE=2           
+RC=250.75)

*lpnp prerad off ctp 3b
.model QLPMOD PNP (             
+IS=7.40964E-16
+BF=90.9
+NF=0.99         
+VAF=36.3423711
+IKF=1.30957E-4  
+NK=0.52
+ISE=6E-16
+NE=1.27089 
+BR=0.697 
+NR=2
+VAR=100  
+IKR=0.1 
+ISC=1E-17
+ NC=2    
+RB=758.578   
+IRB=3.6E-5
+ RBM=100    
+RE=4.096  
+RC=1)

*JFET
.model NJF_TYP NJF (
+ VTO = -1.0    BETA = 6.2E-4   LAMBDA = 0.003 
+ RD = 0.01      RS = 1e-4 
+ CGS = 3E-12    CGD=1.5E-12     IS=5E-10)

.model DMODPNP D (IS = 1.727928319301976e-13
+ N = 1.273993270882892)

.model DMODNPN D (IS = 4.940948456720263e-13
+ N = 1.736958509626848)

*end of the netlist
.end