Title: LM741 /Slewrate / SupplyCurrent (A)
********************************

*Input Voltage Source
*********************
VCC 6 0 DC 15V
VEE 7 0 DC -15V
Vin 1 0 PULSE(0 1 5u 100p 100p 30u 60u)
*********************
*Subcircuit
*X1 26 22 27 28 25
X1 6 7 1 3 3 LM741

*Input
********
.tran 1u 60u
.options timeint method=gear

*Output
.print tran format=noindex file={output_filename}
+ V(1)
+ V(3)
+ I(VEE)
