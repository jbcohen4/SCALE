*Subcircuit name: LM111 Vcc Vee NonInvInput InvInput Output
**************************
.subckt LM111 8 28 35 36 33



*Current source: I<name> <+ node> <- node> [[DC] <value>]
IS1 8 18 10uA

*Resistance: R<name> <+ node> <- node> [model name] <value>
R1 8 6 1400 
R2 8 7 1400
R3 7 9 300
R4 6 9 300
R5 37 5 300
R6 5 10 3400
R7 5 11 3400
R8 8 12 920
R9 8 14 920
R10 30 31 4000
R11 31 32 160
R12 32 34 630
R13 34 0 6
R14 21 28 5100
R15a 21 22 740
R15b 21 26 830
R16 17 22 870
R17 22 23 200
R18 24 28 270
R19 25 28 590
R20 12 15 4000
R21 26 27 970
R22 16 18 270

*Diode: D<name> <anode node (+)> <cathode node (-)> <model name> [area value]
**********************************
*PNP
D1 1 35 DMODSPMOD 1.57 temp=25
D2 2 36 DMODSPMOD 1.54 temp=25
D5a 7 5 DMODPNP 1.3 temp=25
D5b 6 5 DMODPNP 1.3 temp=25
D7 9 14 DMODPNP 0.8 temp=25
D11 14 15 DMODPNP 1.5 temp=25
D14 29 33 DMODSPMOD 2.3 temp=25

*NPN
D3 1 4 DMODNPN 1.6 temp=25
D4 2 4 DMODNPN 1.7 temp=25
D6 8 37 DMODNPN 1.8 temp=25
D8 10 13 DMODNPN 1.7 temp=25
D9 11 13 DMODNPN 1.7 temp=25
D10 12 15 DMODNPN 4.5 temp=25
D12 30 31 DMODNPN 7.5 temp=25
D13 30 29 DMODNPN 1.8 temp=25
D15 32 34 DMODNPN 206 temp=25
D16 34 0 DMODNPN 1.7 temp=25
D18 18 19 DMODNPN 1.8 temp=25
D19 16 17 DMODNPN 1.7 temp=25
D21 23 24 DMODNPN 1.6 temp=25
D22 26 28 DMODNPN 1.7 temp=25
D23 23 25 DMODNPN 1.8 temp=25
D24 27 28 DMODNPN 1.8 temp=25
D25 19 20 DMODNPN 1.7 temp=25
D26 20 28 DMODNPN 1.7 temp=25

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q1 28 35 1 SPMOD 1 temp=25
Q2 28 36 2 SPMOD 0.96 temp=25
Q5a 2 5 7 LPNP_COMPACT 1.3 temp=25
Q5b 1 5 6 LPNP_COMPACT 1.3 temp=25
Q7 14 14 9 LPNP_COMPACT 0.8 temp=25
Q11 30 15 14 LPNP_COMPACT 1.5 temp=25
Q14 28 33 29 SPMOD 1.85 temp=25

Q3 10 1 4 NPN_COMPACT 1.6 temp=25
Q4 11 2 4 NPN_COMPACT 1.7 temp=25
Q6 8 8 37 NPN_COMPACT 1.8 temp=25
Q8 12 10 13 NPN_COMPACT 1.7 temp=25
Q9 14 11 13 NPN_COMPACT 1.7 temp=25
Q10 8 12 15 NPN_COMPACT 4.5 temp=25
Q12 8 30 31 NPN_COMPACT 7.5 temp=25
Q13 30 30 29 NPN_COMPACT 1.8 temp=25
Q15 33 32 34 NPN_COMPACT 206 temp=25
Q16 30 34 0 NPN_COMPACT 1.7 temp=25
Q18 16 18 19 NPN_COMPACT 1.8 temp=25
Q19 15 16 17 NPN_COMPACT 1.7 temp=25
Q21 13 23 24 NPN_COMPACT 1.6 temp=25
Q22 23 26 28 NPN_COMPACT 1.7 temp=25
Q23 4 23 25 NPN_COMPACT 1.8 temp=25
Q24 27 27 28 NPN_COMPACT 1.8 temp=25
Q25 19 19 20 NPN_COMPACT 1.7 temp=25
Q26 20 20 28 NPN_COMPACT 1.7 temp=25

*end of the subcircuit 
.ends


*Library
* npn prerad off ctp 3b
.MODEL  NPN_COMPACT NPN(               
+IS=2.354912E-16
+BF=84.058
+NF=0.986787     
+VAF=351.9861415
+IKF=9.86E-3
+NK=0.47574  
+ISE=7.1029E-15
+NE=2.06453  
+BR=0.697       
+NR=2
+VAR=100
+IKR=0.1         
+ISC=1E-17
+NC=2                          
+RB=140.86       
+IRB=1E-3 
+RBM=50                        
+RE=2           
+RC=250.75)

*lpnp prerad off ctp 3b
.MODEL LPNP_COMPACT PNP (
+IS=7.40964E-16
+BF=90.9
+NF=0.99         
+VAF=36.3423711
+IKF=1.30957E-4  
+NK=0.52
+ISE=6E-16
+NE=1.27089 
+BR=0.697 
+NR=2
+VAR=100  
+IKR=0.1 
+ISC=1E-17
+ NC=2    
+RB=758.578   
+IRB=3.6E-5
+ RBM=100    
+RE=4.096  
+RC=1)

* Substrate PNP
.model SPMOD PNP(
+ IS=1.55E-15
+ BF=1000
+ NF=0.99
+ VAF=36.3423711
+ IKF=7E-5
+ NK=0.52
+ ISE=0.01E-15 
+ NE=1.22
+ BR=0.697
+ NR=2
+ VAR=100
+ IKR=0.1
+ ISC=1E-17
+ NC=2
+ RB=4000 
+ IRB=3.6E-5
+ RBM=100
+ RE=4
+ RC=1)

.model DMODPNP D (IS = {PNP_IS}
+ N = {PNP_N})

.model DMODNPN D (IS = {NPN_IS}
+ N = {NPN_N})

.model DMODSPMOD D (IS = {PNP_IS}
+ N = {PNP_N})

*end of the netlist
.end