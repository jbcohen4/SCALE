*Subcircuit VCC VEE VIN+ VIN- VOUT
**********************************
.subckt LM124_sc 18 8 1 2 15

*Diode: D<name> <anode node (+)> <cathode node (-)> <model name> [area value]
*****************************************************************************

*Current source: I<name> <+ node> <- node> [[DC] <value>]
IS1 19 8 50uA

*PNP
D21         14 7  DMODPNP1 2.12
D51         10 6  DMODPNP1 0.82
D71         11 13  DMODPNP1 0.91
D111        15 9  DMODPNP1 8.51
D15a1       18 19  DMODPNP1 0.87
D15b1       18 19  DMODPNP1 3.22
D16a1       18 19  DMODPNP1 0.29
D16b1       18 19  DMODPNP1 0.29
D171        4 2  DMODPNP1 0.95
D181        5 4  DMODPNP1 0.95
D19a1       18 19  DMODPNP1 0.20
D19b1       18 19  DMODPNP1 0.20
D19c1       18 19  DMODPNP1 0.20
D19d1       18 19  DMODPNP1 0.20
D19e1       18 19  DMODPNP1 0.20
D201       5 3  DMODPNP1 0.99
D211        3 1  DMODPNP1 0.95

D22         14 7  DMODPNP2 2.12
D52         10 6  DMODPNP2 0.82
D72         11 13  DMODPNP2 0.91
D112        15 9  DMODPNP2 8.51
D15a2       18 19  DMODPNP2 0.87
D15b2       18 19  DMODPNP2 3.22
D16a2       18 19  DMODPNP2 0.29
D16b2       18 19  DMODPNP2 0.29
D172       4 2  DMODPNP2 0.95
D182        5 4  DMODPNP2 0.95
D19a2       18 19  DMODPNP2 0.20
D19b2       18 19  DMODPNP2 0.20
D19c2       18 19  DMODPNP2 0.20
D19d2       18 19  DMODPNP2 0.20
D19e2       18 19  DMODPNP2 0.20
D202        5 3  DMODPNP2 0.99
D212        3 1  DMODPNP2 0.95

*NPN
D31         7 8  DMODNPN1 0.48
D41         7 8  DMODNPN1 0.48
D61         10 12  DMODNPN1 0.44
D81         13 8  DMODNPN1 0.54
D91         12 8  DMODNPN1 3.06
D101        13 8  DMODNPN1 1.89
D121        16 15  DMODNPN1 1.44
D131        17 16  DMODNPN1 13.23
D141        9 17  DMODNPN1 1.20

D32         7 8  DMODNPN2 0.48
D42         7 8  DMODNPN2 0.48
D62         10 12  DMODNPN2 0.44
D82         13 8  DMODNPN2 0.54
D92         12 8  DMODNPN2 3.06
D102        13 8  DMODNPN2 1.89
D122        16 15  DMODNPN2 1.44
D132        17 16  DMODNPN2 13.23
D142        9 17  DMODNPN2 1.20

*BJT: Q<name> <collector> <base> <emitter> [substrate] <model name> [area value]
Q2         8 7 14 SPMOD 0.18
Q3         7 7 8 NPN_compact 0.48
Q4         6 7 8 NPN_compact 0.48
Q5         8 6 10 SPMOD 0.03
Q6         11 10 12 NPN_compact 0.44
Q7         8 13 11 SPMOD 0.03
Q8         13 13 8 NPN_compact 0.54
Q9         9 12 8 NPN_compact 3.06
Q10        15 13 8 NPN_compact 1.89
Q11        8 9 15 SPMOD 1.04
Q12        9 16 15 NPN_compact 1.44
Q13        18 17 16 NPN_compact 13.23
Q14        18 9 17 NPN_compact 1.20
Q15a       19 19 18 LPNP_compact 0.87
Q15b       9 19 18 LPNP_compact 3.22
Q16a       13 19 18 LPNP_compact 0.29

Q16b       11 19 18 LPNP_compact 0.29
Q17        8 2 4 SPMOD 0.04
Q18        7 4 5 LPNP_compact 0.95
Q19a       5 19 18 LPNP_compact 0.20
Q19b       3 19 18 LPNP_compact 0.20
Q19c       4 19 18 LPNP_compact 0.20
Q19d       14 19 18 LPNP_compact 0.20
Q19e       10 19 18 LPNP_compact 0.20
Q20        6 3 5 LPNP_compact 0.99
Q21        8 1 3 SPMOD 0.04

*Resistance: R<name> <+ node> <- node> [model name] <value>
R1          17 16 40K
R2          16 15 25

*Capacitance: C<name> <+ node> <- node> [model name] <value> + [IC=<initial value>]
C1 9 6 18p

.ends LM124_sc

.model NPN_COMPACT NPN(               
+IS=2.354912E-16
+BF=84.058
+NF=0.986787     
+VAF=351.9861415
+IKF=9.86E-3
+NK=0.47574  
+ISE=7.1029E-15
+NE=2.06453  
+BR=0.697       
+NR=2
+VAR=100
+IKR=0.1         
+ISC=1E-17
+NC=2                          
+RB=140.86       
+IRB=1E-3 
+RBM=50                        
+RE=2           
+RC=250.75)

.model LPNP_compact PNP (
+IS=7.40964E-16
+BF=90.9
+NF=0.99         
+VAF=36.3423711
+IKF=1.30957E-4  
+NK=0.52
+ISE=6E-16
+NE=1.27089 
+BR=0.697 
+NR=2
+VAR=100  
+IKR=0.1 
+ISC=1E-17
+ NC=2    
+RB=758.578   
+IRB=3.6E-5
+ RBM=100    
+RE=4.096  
+RC=1)
 
.model SPMOD PNP(
+ IS=11E-15
+ BF=8500
+ NF=0.99
+ VAF=36.3423711
+ IKF=900E-6
+ NK=0.52
+ ISE=0.08E-15 
+ NE=1.3
+ BR=0.697
+ NR=2
+ VAR=100
+ IKR=0.1
+ ISC=1E-17
+ NC=2
+ RB=3058.578 
+ IRB=3.6E-5
+ RBM=100
+ RE=4
+ RC=1)

.model DMODPNP1 D (IS = {PNP_IS_1}
+ N = {PNP_N_1})

.model DMODPNP2 D (IS = {PNP_IS_2}
+ N = {PNP_N_2})

.model DMODNPN1 D (IS = {NPN_IS_1}
+ N = {NPN_N_1})

.model DMODNPN2 D (IS = {NPN_IS_2}
+ N = {NPN_N_2})


*end of the list
.end


